Library IEEE;
use ieee.std_logic_1164.ALL;

Entity my_gates is
	generic (gate_delay : time := 10.0 ns);
	port(a,b: in std_logic;
		o: out std_logic);
end entity;

Architecture xor_arch of my_gates is
	begin 
		o <= a xor b after gate_delay;
	end xor_arch;


Architecture and_arch of my_gates is
	begin
		o <= a and b after gate_delay;
	end and_arch; 

Architecture or_arch of my_gates is
	begin
		o <= a or b after gate_delay;
	end or_arch; 